    Mac OS X            	   2  �     �                                    ATTR��  �   �   I                  �   9  com.apple.quarantine    �     com.apple.lastuseddate#PS 0B-0083;63c8741b;Safari;49E90396-DEC0-450B-A3E8-F491CD73B3A8�l�e    ^Zo'                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          This resource fork intentionally left blank                                                                                                                                                                                                                            ��